
class Generator;

  

endclass


class Generator;

  transaction trans_queue[$];
  
  function new();
  
  endfunction
  
  

endclass


`ifndef CALC_IF_DEFINE
`define CALC_IF_DEFINE








`endif

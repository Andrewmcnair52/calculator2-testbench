
class Generator;

  trans_queue[$];
  
  function new();
  
  endfunction
  
  

endclass
